library ieee;
use ieee.std_logic_1164.all;

package DataStructures is
	type Coordinates is record
		x : integer;
		y : integer;
	end record;

	type ShellObject is record
		cord : Coordinates;
		enabled : std_logic;
	end record;


	type ArrayOfShells is array(0 to 9) of ShellObject;

	type ShipType is record
		color : std_logic_vector (23 downto 0);
		value : integer;

		ship_image_width : integer;
		ship_image_height : integer;
	end record;

	type ShipObject is record
		pos1 : Coordinates;
		ship_type : ShipType;
	end record;

	type ShipArray is array(0 to 4) of ShipObject;

	constant destroyer : ShipType := (
		color => "011111000000000000011111",
		value => 1,
		ship_image_width => 11,
		ship_image_height => 114
	);
	constant battleShip : ShipType := (
		color => "000000011111000000011111",
		value => 5,
		ship_image_width => 20,
		ship_image_height => 65
	);
	constant civilShip : ShipType := (
		color => "000000000000001111111111",
		value => - 2,
		ship_image_width => 20,
		ship_image_height => 65
	);

	type GraphicMemoryType is array(0 to 1300) of std_logic_vector(7 downto 0);
end package DataStructures;



package body DataStructures is
end package body DataStructures;